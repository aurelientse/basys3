//------------------------------------------------------
//------------------------------------------------------
// FILENAME : parameters.svh
// TESTBENCH PARAMETER FOR BLINK LED 
//-----------------------------------------------------
//-----------------------------------------------------

`define PERIOD 10  // 100MHz (Basys3 clock frequency)